/*
*  File            :   avalon_drv.sv
*  Autor           :   Vlasov D.V.
*  Data            :   2020.01.09
*  Language        :   SystemVerilog
*  Description     :   This is avalon interface driver 
*  Copyright(c)    :   2019 - 2020 Vlasov D.V.
*/

`ifndef AVALON_DRV__SV
`define AVALON_DRV__SV

class avalon_drv extends dvv_drv #(ctrl_trans);
    `OBJ_BEGIN( avalon_drv )

    virtual avalon_if           vif;

    ctrl_trans                  item;

    avalon_mth                  mth;

    dvv_aep #(logic [15 : 0])   u_mon_aep;

    uart_struct                 h_uart = new_uart( 0 , 2 );

    extern function new(string name = "", dvv_bc parent = null);

    extern task write_reg(logic [31 : 0] w_addr, logic [31 : 0] w_data);
    extern task read_reg(logic [31 : 0] r_addr, output logic [31 : 0] r_data);

    extern task build();
    extern task run();
    
endclass : avalon_drv

function avalon_drv::new(string name = "", dvv_bc parent = null);
    super.new(name,parent);
    u_mon_aep = new();
endfunction : new

task avalon_drv::build();
    if( !dvv_res_db#(virtual avalon_if)::get_res_db("avalon_if_0",vif) )
        $fatal();

    mth = avalon_mth::create::create_obj("[ AVALON DRV MTH ]", this);
    mth.vif = vif;

    item = ctrl_trans::create::create_obj("[ AVALON ITEM ]", this);
    item_sock = new();

    $display("%s build complete", this.fname);
endtask : build

task avalon_drv::write_reg(logic [31 : 0] w_addr, logic [31 : 0] w_data);
    mth.set_address(w_addr);
    mth.set_writedata(w_data);
    mth.set_chipselect('1);
    mth.set_write('1);
    mth.wait_clk();
    mth.set_chipselect('0);
    mth.set_write('0);
endtask : write_reg

task avalon_drv::read_reg(logic [31 : 0] r_addr, output logic [31 : 0] r_data);
    mth.set_address(r_addr);
    mth.set_chipselect('1);
    mth.set_write('0);
    mth.wait_clk();
    mth.set_chipselect('0);
    mth.wait_clk();
    mth.set_write('0);
    r_data = mth.get_readdata();
endtask : read_reg

task avalon_drv::run();
    mth.wait_reset();

    h_uart.cr_c.data.rx_fifo_lvl = '0;
    h_uart.cr_c.data.tx_fifo_lvl = '0;
    h_uart.cr_c.data.rec_en      = '0;
    h_uart.cr_c.data.tr_en       = '1;

    write_reg(h_uart.cr_c.addr, h_uart.cr_c.data);

    item_sock.trig_sock();
    forever
    begin
        item_sock.rec_msg(item);
        
        h_uart.tx_rx_c.data = item.data;
        h_uart.dfr_c.data = item.freq;

        write_reg(h_uart.dfr_c.addr, h_uart.dfr_c.data);

        u_mon_aep.write(h_uart.dfr_c.data);
        
        write_reg(h_uart.tx_rx_c.addr, h_uart.tx_rx_c.data);

        for(;;)
        begin
            read_reg(h_uart.cr_c.addr, h_uart.cr_c.data);
            if( h_uart.cr_c.data.tx_full == 0 )
                break;
        end

        item_sock.trig_sock();
    end
endtask : run

`endif // AVALON_DRV__SV
